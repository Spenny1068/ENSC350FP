library ieee;
Use ieee.std_logic_1164.all;

Entity LogicUnit is
Generic ( N : natural := 64);
Port(A, B: in std_logic_vector(N-1 downto 0);
	Y: out std_logic_vector(N-1 downto 0);
	LogicFN: in std_logic_vector(1 downto 0));
End Entity LogicUnit;

Architecture rtl of LogicUnit is
	Signal PassB, AxorB, AorB, AandB : std_logic_vector(N-1 downto 0);
Begin

gen: 	for i in N-1 downto 0 generate
	PassB(i) <= B(i);
	AxorB(i) <= A(i) XOR B(i);
	AorB(i) <= A(i) OR B(i);
	AandB(i) <= A(i) AND B(i);
	end generate gen;
	
	with LogicFN select
	Y <= PassB when "00", AxorB when "01", AorB when "10", AandB when others;

End Architecture rtl;